/**********************************************************************************
* * Módulo: main
*
* Descrição: 
* Este é o módulo de topo que integra um sistema de processamento de imagens 
* em uma FPGA. Ele gerencia a leitura de uma imagem de uma ROM, o envio para 
* um coprocessador que aplica algoritmos de redimensionamento (zoom in/out) 
* selecionados por chaves (SW), o armazenamento da imagem processada em uma RAM
* e, por fim, a exibição do resultado em um monitor VGA. O módulo também 
* controla a geração de clocks e a lógica de reset automático baseada nas chaves.
* O processamento inicia automaticamente ao selecionar um algoritmo nas chaves SW.
*
**********************************************************************************/
module main (
    input  wire [9:2] SW,
    input  wire [1:0] boton, // Botão ainda presente na interface, mas boton[0] não é usado para start
    input  wire clk_50,
    output wire [9:0] LEDR,
    output wire hsync,
    output wire vsync,
    output wire [7:0] red,
    output wire [7:0] green,
    output wire [7:0] blue,
    output wire sync,
    output wire clk,
    output wire blank
);

    assign LEDR = SW;
    reg clk_25_reg = 0;
    
    always @(posedge clk_50) begin
        clk_25_reg <= ~clk_25_reg;
    end
    
    // --- Lógica de Reset Automático ao Mudar as Chaves ---
    reg [7:0] sw_prev = 0;         
    reg       auto_reset_flag = 0; 
    reg [3:0] reset_counter = 0;   
    
    wire sw_changed = (sw_prev != SW[8:2]);
    
    always @(posedge clk_25_reg) begin
        sw_prev <= SW[8:2]; 
        
        if (sw_changed) begin
            auto_reset_flag <= 1'b1;     
            reset_counter <= 4'd15;      
        end else if (reset_counter > 0) begin
            reset_counter <= reset_counter - 1;
            if (reset_counter == 1)
                auto_reset_flag <= 1'b0; 
        end
    end
    
    wire reset = SW[9] || auto_reset_flag;
    
    // --- PLL ---
    wire clock_100; 
    wire locked; 
    pll100_0002 pll100_inst (
        .refclk   (clk_50),    
        .rst      (1'b0), // Idealmente, conectar ao reset do sistema se necessário
        .outclk_0 (clock_100), 
        .locked   (locked)     
    );

    // --- Sinais VGA ---
    wire [10:0] next_x;
    wire [10:0] next_y;
    reg [10:0] x_delayed;
    reg [10:0] y_delayed;

    always @(posedge clk_25_reg) begin
        x_delayed <= next_x;
        y_delayed <= next_y;
    end
    
    // --- Constantes ---
    localparam IMG_WIDTH_PEQ8  = 20;
    localparam IMG_HEIGHT_PEQ8 = 15;
    localparam IMG_WIDTH_PEQ4  = 40;
    localparam IMG_HEIGHT_PEQ4 = 30;
    localparam IMG_WIDTH_PEQ   = 80;
    localparam IMG_HEIGHT_PEQ  = 60;
    localparam IMG_WIDTH_OR    = 160;
    localparam IMG_HEIGHT_OR   = 120;
    localparam IMG_WIDTH_GRA   = 320;
    localparam IMG_HEIGHT_GRA  = 240;      
    localparam IMG_WIDTH_GRA4  = 640;
    localparam IMG_HEIGHT_GRA4 = 480;
    localparam IMG_TOTAL_PIXELS_OR = IMG_WIDTH_OR * IMG_HEIGHT_OR;

    // --- Sinais Coprocessador ---
    wire        processing_done;
    wire        coproc_pixel_in_ready;
    
    wire modo_processamento_ativo = (SW[5:2] != 4'b0000); // Modo ativo se alguma chave de algoritmo estiver ligada

    // --- Contador de Leitura da ROM (agora inicia com modo_processamento_ativo) ---
    reg [18:0] rom_addr_counter = 0;
    always @(posedge clk_25_reg or posedge reset) begin
        if (reset) begin
            rom_addr_counter <= 0;
        // MODIFICADO: Remove 'boton[0]', adiciona 'modo_processamento_ativo'
        end else if (modo_processamento_ativo && !processing_done && rom_addr_counter < IMG_TOTAL_PIXELS_OR && coproc_pixel_in_ready) begin
            rom_addr_counter <= rom_addr_counter + 1;
        end
        // O contador para automaticamente quando as condições não são mais atendidas ou reseta com 'reset'
    end

    // --- Lógica de Endereçamento VGA ---
    reg [18:0] ram_address_read;
    // ... (definições de dentro_img_xxx e ram_addr_xxx permanecem iguais) ...
    wire dentro_img_peq = (x_delayed < IMG_WIDTH_PEQ) && (y_delayed < IMG_HEIGHT_PEQ);
    wire [18:0] ram_addr_peq = dentro_img_peq ? (y_delayed * IMG_WIDTH_PEQ + x_delayed) : 19'd0;
    wire dentro_img_peq4 = (x_delayed < IMG_WIDTH_PEQ4) && (y_delayed < IMG_HEIGHT_PEQ4);
    wire [18:0] ram_addr_peq4 = dentro_img_peq4 ? (y_delayed * IMG_WIDTH_PEQ4 + x_delayed) : 19'd0;
    wire dentro_img_peq8 = (x_delayed < IMG_WIDTH_PEQ8) && (y_delayed < IMG_HEIGHT_PEQ8);
    wire [18:0] ram_addr_peq8 = dentro_img_peq8 ? (y_delayed * IMG_WIDTH_PEQ8 + x_delayed) : 19'd0;
    wire dentro_img_or_display = (x_delayed < IMG_WIDTH_OR) && (y_delayed < IMG_HEIGHT_OR);
    wire [18:0] ram_addr_or = dentro_img_or_display ? (y_delayed * IMG_WIDTH_OR + x_delayed) : 19'd0;
    wire dentro_img_gra = (x_delayed < IMG_WIDTH_GRA) && (y_delayed < IMG_HEIGHT_GRA);
    wire [18:0] ram_addr_gra = dentro_img_gra ? (y_delayed * IMG_WIDTH_GRA + x_delayed) : 19'd0;
    wire dentro_img_gra4 = (x_delayed < IMG_WIDTH_GRA4) && (y_delayed < IMG_HEIGHT_GRA4);
    wire [18:0] ram_addr_gra4 = dentro_img_gra4 ? (y_delayed * IMG_WIDTH_GRA4 + x_delayed) : 19'd0;
    
    always @(*) begin
        // Define um valor padrão para evitar latches
        ram_address_read = ram_addr_or; 
    
        case (SW[8:7]) 
            2'b01: begin 
                case (SW[5:2])
                    4'b0001:  ram_address_read = ram_addr_gra4;
                    default:  ram_address_read = ram_addr_or;
                endcase
            end
            
            2'b10: begin 
                case (SW[5:2])
                    4'b0001:  ram_address_read = ram_addr_gra4; 
                    default:  ram_address_read = ram_addr_or;
                endcase
            end
            
            default: begin 
                case (SW[5:2])
                    4'b0001, 4'b0010:  ram_address_read = ram_addr_gra;
                    4'b0100, 4'b1000:  ram_address_read = ram_addr_peq;
                    default:           ram_address_read = ram_addr_or;
                endcase
            end
        endcase
    end
    
    // --- Lógica de Seleção de Fonte de Dados ---
    wire [7:0] saida_rom;
    wire [18:0] address_rom;
    wire [7:0]  entrada_vga;
    reg  process_done_latch = 0; // Latch para indicar que o processamento terminou

    assign address_rom = modo_processamento_ativo ? rom_addr_counter : ram_addr_or;
    assign entrada_vga = (modo_processamento_ativo && process_done_latch) ? ram_q : saida_rom;
    
    // --- Instância da ROM ---
    imagem rom_inst_OR (
        .address(address_rom),
        .clock(clock_100),
        .q(saida_rom)
    );

    // --- Instância do Coprocessador (agora 'start' depende do modo) ---
    wire [7:0] pixel_coproc_out;
    wire       pixel_coproc_valid;
    
    // MODIFICADO: Sinal 'start' agora é ativado pelo modo e enquanto não terminou
    wire coproc_start_signal = modo_processamento_ativo && !process_done_latch; 
    
    coprocessador coprocessador_inst (
        .clk(clk_25_reg), 
        .resetn(~reset), 
        .start(coproc_start_signal), // Conecta o novo sinal de start
        .largura_in(IMG_WIDTH_OR),
        .altura_in(IMG_HEIGHT_OR), 
        .SW(SW[5:2]), 
        .escala(SW[8:7]),
        .pixel_in(saida_rom),
        .pixel_out(pixel_coproc_out), 
        .pixel_out_valid(pixel_coproc_valid),
        .processing_done(processing_done), 
        .pixel_in_ready(coproc_pixel_in_ready)
    );

    // --- Controle da RAM de Saída ---
    reg  [18:0] pixel_write_count = 0;
    
    always @(posedge clk_25_reg or posedge reset) begin
        if (reset) begin
            pixel_write_count  <= 0;
            process_done_latch <= 0;
        end else begin
            // Só escreve na RAM se o coprocessador fornecer um pixel válido E o processamento não tiver terminado
            if (pixel_coproc_valid && !process_done_latch) begin
                pixel_write_count <= pixel_write_count + 1;
            end
            // Trava o sinal de 'done' quando o coprocessador indicar que terminou
            if (processing_done) begin
                process_done_latch <= 1'b1; 
            end
        end
    end

    wire [18:0] ram_address_write = pixel_write_count;
    // O endereço para a RAM alterna entre escrita (durante proc.) e leitura (após proc.)
    wire [18:0] ram_address = process_done_latch ? ram_address_read : ram_address_write; 
    // Habilita escrita na RAM apenas durante o processamento e quando há pixel válido
    wire        escrita     = pixel_coproc_valid && !process_done_latch; 
    wire [7:0]  ram_q;
    
    // --- Instância da RAM ---
    ram_pri ram_inst (
        .address(ram_address),
        .clock(clock_100), // Usando clock rápido para a RAM
        .data(pixel_coproc_out),   
        .wren(escrita), 
        .q(ram_q)
    );

    // --- Instância do VGA ---
    vga_module vga_inst (
        .clock(clk_25_reg), 
        .reset(reset), 
        .color_in(entrada_vga), // A fonte já foi selecionada corretamente acima
        .next_x(next_x),
        .next_y(next_y), 
        .hsync(hsync), 
        .vsync(vsync), 
        .red(red), 
        .green(green),
        .blue(blue), 
        .sync(sync), 
        .clk(clk), 
        .blank(blank)
    );

endmodule